module part1 (input Clock, input Enable, input Reset, output [7:0] CounterValue);
