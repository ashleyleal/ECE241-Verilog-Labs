module part3(clock, reset, ParallelLoadn, RotateRight, ASRight, Data IN, Q);


